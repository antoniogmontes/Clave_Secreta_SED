--LAURA BUTANERA